library verilog;
use verilog.vl_types.all;
entity control_module_tb is
end control_module_tb;
