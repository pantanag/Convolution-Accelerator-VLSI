library verilog;
use verilog.vl_types.all;
entity convolution_module_tb is
end convolution_module_tb;
